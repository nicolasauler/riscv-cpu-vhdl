library ieee;
use ieee.std_logic_1164.all;
use std.textio.all;
use ieee.numeric_std.all;
use ieee.std_logic_textio.all;

entity instrmem is 
    port(
        a:      in  std_logic_vector(31 downto 0);
        rd:     out std_logic_vector(31 downto 0)
    );
end entity instrmem;

architecture behavioural of instrmem is 

type ramtype is array (63 downto 0) of std_logic_vector(31 downto 0);

constant mem: ramtype := (
0   => "00000000000000000010000010000011", -- lw x1, 0(x0) -> carrega 7
1   => "00000000000000001000000100110011", -- add x2, x1, x0 -> x2 = 7
2   => "00000000000000001000000110110011", -- add x3, x1, x0 -> x3 = 7
3   => "01000000000100010000000110110011", -- sub x3, x2, x1 -> x3 = 0
4   => "00000000000100010111000010110011", -- and x1, x2, x1 -> x1 = x1
5   => "00000000000000110000100110001111", -- beq x3, x0, 8
6   => "00000000001000001000000010110011", -- add x1, x1, x2 -> x1 = 14
7   => "00000010000100000010010000100011", -- sw x1, 40(x0) -> if branch, x1 = 7, else x1=14
8   => "00000000010000100000000110001111", -- beq x2, x2, 0
9   => "00000000000000000000000000000000", -- 
10  => "00000000000000000000000000000000", -- 
11  => "00000000000000000000000000000000", -- 
12  => "00000000000000000000000000000000",
13  => "00000000000000000000000000000000",
14  => "00000000000000000000000000000000",
15  => "00000000000000000000000000000000",
16  => "00000000000000000000000000000000",
17  => "00000000000000000000000000000000",
18  => "00000000000000000000000000000000",
19  => "00000000000000000000000000000000",
20  => "00000000000000000000000000000000",
21  => "00000000000000000000000000000000",
22  => "00000000000000000000000000000000",
23  => "00000000000000000000000000000000",
24  => "00000000000000000000000000000000",
25  => "00000000000000000000000000000000",
26  => "00000000000000000000000000000000",
27  => "00000000000000000000000000000000",
28  => "00000000000000000000000000000000",
29  => "00000000000000000000000000000000",
30  => "00000000000000000000000000000000",
31  => "00000000000000000000000000000000",
32  => "00000000000000000000000000000000",
33  => "00000000000000000000000000000000",
34  => "00000000000000000000000000000000",
35  => "00000000000000000000000000000000",
36  => "00000000000000000000000000000000",
37  => "00000000000000000000000000000000",
38  => "00000000000000000000000000000000",
39  => "00000000000000000000000000000000",
40  => "00000000000000000000000000000000",
41  => "00000000000000000000000000000000",
42  => "00000000000000000000000000000000",
43  => "00000000000000000000000000000000",
44  => "00000000000000000000000000000000",
45  => "00000000000000000000000000000000",
46  => "00000000000000000000000000000000",
47  => "00000000000000000000000000000000",
48  => "00000000000000000000000000000000",
49  => "00000000000000000000000000000000",
50  => "00000000000000000000000000000000",
51  => "00000000000000000000000000000000",
52  => "00000000000000000000000000000000",
53  => "00000000000000000000000000000000",
54  => "00000000000000000000000000000000",
55  => "00000000000000000000000000000000",
56  => "00000000000000000000000000000000",
57  => "00000000000000000000000000000000",
58  => "00000000000000000000000000000000",
59  => "00000000000000000000000000000000",
60  => "00000000000000000000000000000000",
61  => "00000000000000000000000000000000",
62  => "00000000000000000000000000000000",
63  => "00000000000000000000000000000000"
);

begin

    -- read memory
    process(a)
    begin
        rd <= mem(to_integer(unsigned(a(31 downto 2))));
    end process;

end architecture behavioural;
